--Author : Abel DIDOUH
--Schema 2
---------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
---------------------------------------------------------------------------------------------------
entity ctr_tempo_entity is 
    generic(
        X : 
    )