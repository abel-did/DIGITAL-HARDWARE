    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.apple.TextEncoding      �     com.apple.lastuseddate#PS    UTF-8;134217984��'d    ��.    